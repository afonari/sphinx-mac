netcdf keyword3 {
variables:
	real f ;
	long l ;
}
